/**
 * Copyright (c) 2016 C. Brett Witherspoon
 */
package funct3;

    localparam BEQ   = 3'b000;
    localparam LB    = 3'b000;
    localparam SB    = 3'b000;
    localparam ADD   = 3'b000;
    localparam SUB   = 3'b000;
    localparam BNE   = 3'b001;
    localparam LH    = 3'b001;
    localparam SH    = 3'b001;
    localparam SLL   = 3'b001;
    localparam LW    = 3'b010;
    localparam SW    = 3'b010;
    localparam SLT   = 3'b010;
    localparam SLTU  = 3'b011;
    localparam SLTIU = 3'b011;
    localparam BLT   = 3'b100;
    localparam XOR   = 3'b100;
    localparam LBU   = 3'b100;
    localparam BGE   = 3'b101;
    localparam LHU   = 3'b101;
    localparam SRL   = 3'b101;
    localparam SRA   = 3'b101;
    localparam BLTU  = 3'b110;
    localparam OR    = 3'b110;
    localparam BGEU  = 3'b111;
    localparam AND   = 3'b111;

endpackage
