/**
 * Module: writeback
 */
module writeback;


endmodule
