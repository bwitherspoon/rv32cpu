/**
 * Module: core
 * 
 * The processor core.
 */
module core (
    input logic clk,
    input logic resetn
);

endmodule


