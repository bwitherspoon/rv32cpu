/**
 * Package: riscv
 */
package riscv;

    localparam WORD_WIDTH = 32;
    localparam REGS_ADDR_WIDTH = 5;
    localparam REGS_DATA_WIDTH = WORD_WIDTH;
    localparam IMEM_ADDR_WIDTH = 9;
    localparam IMEM_DATA_WIDTH = WORD_WIDTH;
    
endpackage


