/**
 * Package: funct7
 */
package funct7;

    typedef logic [6:0] funct7_t;
    
    localparam funct7_t ADDSRL = 'b000000;
    localparam funct7_t SUBSRA = 'b010000;
    localparam funct7_t MULDIV = 'b000001;

endpackage


